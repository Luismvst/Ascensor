Multiplexor.vhd

entity Multiplex is
port (
	accion_motor: in std_logic;
	accio)