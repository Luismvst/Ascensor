Display7seg.vhd

--Lo haremos al final